library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ctrlUnit is
    port (
        instr : in unsigned (15 downto 0) := "0000000000000000";
        ULAop : out unsigned (1 downto 0) := "00" -- selecao de operacoes da ULA
        ULA_srcA : out std_logic := '0'; -- MUX source do RegA da ULA
        ULA_srcB : out std_logic := '0'; -- MUX source do RegB da ULA
        regWr_en : out std_logic := '0'; -- wr_en do regBank
        regWr_src : out std_logic := '0'; -- MUX memória ou acumulador
        regWr_address : out std_logic := out unsigned(2 downto 0) -- endereco banco de registradores
        ACM_wr_en : out std_logic := '0'; -- wr_en do ACM
        PC_src : out std_logic := '0'; -- MUX source do PC
        PC_wr_en : out std_logic := '0'; -- wr_en do PC
    );
end entity;

architecture ctrlUnit_Arch of ctrlUnit is

    signal opcode : unsigned(3 downto 0);
    signal funct : std_logic := '0';
    signal ULA_srcA : std_logic := '0';
    signal ULA_op : unsigned(1 downto 0);
begin
    opcode <= instr(15 downto 11);
    funct <= instr(10);
    reg_address <= instr(10 downto 8);

    -- OP_ctrl
    ULA_op <= opcode(1 downto 0); -- instr(12 downto 11)

    -- funct = 1 (com imediato)
    ULA_srcA <= funct;

    -- 1 quando LD para Acumulador ou Mov para Acumulador (Reg ZERO)
    ULA_srcB <= '1' when opcode = "0100" and funct = '1' else
        '1' when opcode = "1100" and funct = '1' else
        '0';

    -- 1 quando LD para Registrador
    regWr_src <= '1' when opcode = "1100" and funct = '0' else
        '0';

    -- 1 quando LD para Registrador e MOV para Registrador
    regWr_en <= '1' when opcode = "0100" and funct = '0' else
        '1' when opcode = "1100" and funct = '0' else
        '0';

    --- 0 quando CMP, LD para Registrador, MOV para Registrador e JMP
    ACM_wr_en <= '0' when opcode = "0001" and funct = '0' else
        '0' when opcode = "0100" and funct = '0' else
        '0' when opcode = "1100" and funct = '0' else
        '0' when opcode = "1111" else
        '1';

    -- Sempre, por enquanto
    PC_wr_en <= '1';

    -- 1 quando JMP
    PC_src <= '1' when opcode = "1111" else
    '0';

end architecture;